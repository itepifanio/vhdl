-- Aula 04 - exercicio 1
--package exercicio_1 is
--	type BYTE is array(3 downto 0) of BIT;
--end exercicio_1;

entity exercicio_1 is 
end exercicio_1;

architecture Behavior of exercicio_1 is 
begin
end Behavior;