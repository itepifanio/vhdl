-- Por estar utilizando o EDA playground não consegui rodar as simulações, isso será feito posteriormente
